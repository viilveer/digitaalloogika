library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity JUHTAUTOMAAT is 
    Port ( -- sisendid siia
    	); --4 bit output 
end JUHTAUTOMAAT;

architecture toplevel of JUHTAUTOMAAT is
-- sisendsignaalid siia

-- komponendid siia 
begin --beginning of the architecture

-- port maps here
	
end toplevel;